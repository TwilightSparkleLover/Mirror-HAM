[Font]
Font=
Name=Courier New
Size=9
[Assembler]
Assembler=
ForeGround=$800000
BackGround=$FFFFFF
[Comment]
Comment=
ForeGround=$008000
BackGround=$FFFFFF
[Directive]
Directive=
ForeGround=$FF0000
BackGround=$FFFFFF
[Identifier]
Identifier=
ForeGround=$000000
BackGround=$FFFFFF
[Invalid]
Invalid=
ForeGround=$000000
BackGround=$FFFFFF
[Key]
Key=
ForeGround=$FF0000
BackGround=$FFFFFF
[Number]
Number=
ForeGround=$0000FF
BackGround=$FFFFFF
[Space]
Space=
ForeGround=$FFFFFF
BackGround=$FFFFFF
[String]
String=
ForeGround=$808080
BackGround=$FFFFFF
[Symbol]
Symbol=
ForeGround=$000000
BackGround=$FFFFFF
[Editor]
Editor=
ForeGround=$000000
BackGround=$FFFFFF
