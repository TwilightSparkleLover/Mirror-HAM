[Font]
Name=Courier New
Size=9

[Assembler]
ForeGround=$00ff00
BackGround=$000000

[Comment]
ForeGround=$c0c0c0
BackGround=$000000

[Directive]
ForeGround=$ffff00
BackGround=$000000

[Identifier]
ForeGround=$80000005
BackGround=$000000

[Invalid]
ForeGround=$ffffff
BackGround=$FF0000

[Key]
ForeGround=$ffff00
BackGround=$000000

[Number]
ForeGround=$ff00ff
BackGround=$000000

[Space]
ForeGround=$000000
BackGround=$000000

[String]
ForeGround=$00ffff
BackGround=$000000

[Symbol]
ForeGround=$ffff00
BackGround=$000000

[Editor]
ForeGround=$000000
BackGround=$000000