[Font]
Font=
Name=Courier New
Size=9

[Assembler]
Assembler=
ForeGround=$000000
BackGround=$FFFFFF

[Comment]
Comment=
ForeGround=$800000
BackGround=$FFFFFF

[Directive]
Directive=
ForeGround=$000000
BackGround=$FFFFFF

[Identifier]
Identifier=
ForeGround=$000000
BackGround=$FFFFFF

[Invalid]
Invalid=
ForeGround=$FFFFFF
BackGround=$0000FF

[Key]
Key=
ForeGround=$000000
BackGround=$FFFFFF

[Number]
Number=
ForeGround=$800000
BackGround=$FFFFFF

[Space]
Space=
ForeGround=$FFFFFF
BackGround=$FFFFFF

[String]
String=
ForeGround=$800000
BackGround=$FFFFFF

[Symbol]
Symbol=
ForeGround=$000000
BackGround=$FFFFFF

[Editor]
Editor=
ForeGround=$000000
BackGround=$FFFFFF
